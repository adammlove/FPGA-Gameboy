module inputs(
input wire [7:0] button
);

endmodule