module PPU();

endmodule